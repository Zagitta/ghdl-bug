library ieee;
use ieee.std_logic_1164.all;

library work;
use work.pkg1.all;
use work.pkg2.all;

entity top is
port (
    clk : in std_logic
);
end top;

architecture arch of top is
begin
end architecture;
