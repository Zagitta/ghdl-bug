package pkg2 is

end pkg2;
