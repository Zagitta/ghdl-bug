package pkg1 is
end pkg1;
